library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity something is
    port(
        signal1     : in    std_logic;
        signal2     : out   std_logic
    );
end something;

architecture rtl of something is

    #Constants
    #signals

begin





end something;
